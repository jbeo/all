
library IEEE;

